/**
 * testbench template
 *
 * @version: 0.1
 * @author : Gabriel Villanova N. M.
 */

 module tb;

  // main block
  initial begin
    $display("\n\nWhat do wanna test?\n");
    $finish();
  end

endmodule