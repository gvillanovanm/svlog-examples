/**
 * testbench template
 *
 * @version: 0.1
 * @author : Gabriel Villanova N. M.
 */
module tb;
    import uvm_pkg::*;
    `include "uvm_macros.svh"  

    import eg_pkg::*;

    initial begin
        run_test();
    end
endmodule