package eg_pkg;
  // uvm
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  // eg
  `include "eg_seq_item.svh"
  `include "eg_sequence.svh"
  `include "eg_source.svh"
  `include "eg_sink.svh"
  `include "eg_env.svh"
  `include "eg_test_basic.svh"

endpackage
