/**
 * DUT template
 *
 * @version: 0.1
 * @author : Gabriel Villanova N. M.
 */

module dut #(
  // parameters
) (
  // port_list
);
  
endmodule